`ifndef SPMV_MACROS
`define SPMV_MACROS

// DCP Macros (Assume Fixed to Default)
`define DCP_PADDR_MASK 39:0
`define DCP_NOC_RES_DATA_SIZE 512

`define MAX_DIM_LEN 1024
`define DIM_W       10
`define NNZ_W       20

`endif 